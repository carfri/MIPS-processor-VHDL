library IEEE;
use IEEE.std_logic_1164.all;

entity programmemory is
  port( address:in std_logic_vector(31 downto 0);
        instruction: out std_logic_vector(31 downto 0)
        );
end programmemory;

architecture behav of programmemory is
begin

with address select
  instruction <=
		--	"00100000001000001111111111111000" when X"00000000",  --addi r0,r1,-8
       --  "00100000010000010000000000000011" when X"00000004",  --addi r1,r2,3
		 --  "00000000000000010001000000100000" when X"00000008",  --add r2,r0,r1
       --  "00000000001000000001100000100010" when X"0000000c",  --sub r3,r1,r0
		 --  "00000000010000110010000000101010" when X"00000010",  --slt r4,r2,r3
		--	"00101000010001001111111111110111" when X"00000014",  --slti r4,r2,-9
		--	"00000000010000110010000000101010" when X"00000018",  --slt r4,r2,r3
		--	"00000000100001100010100000100101" when X"0000001c",  --or  r5,r4,r6
		--	"00000000101000010011000000100100" when X"00000020",  --and r6,r5,r1
		--	"10101100111000100000000000000000" when X"00000024",  --sw r2,0(r7)
		--	"10001100111010000000000000000000" when X"00000028",	--lw r8,0(r7)
		--	"10101110001000110000000000000100" when X"0000002c",	--sw r3,4(r9)
		--	"10001101010010010000000000000100" when X"00000030",	--lw r9,4(r10) 
			--Muliplication of 5 and 3
		--	"00100000001010100000000000000010" when X"00000034",  --addi r10,r1,2
		--	"00100000001010110000000000000000" when X"00000038",	--addi r11,r1,0
		--	"00100000001011001111111111111101" when X"0000003c",	--addi r12,r1,-3
		--	"00100000001011011111111111111101" when X"00000040",	--addi r13,r1,-3
			
		--	"00010001100010110000000000000011" when X"00000044",	--beq r12, r11,exit
		--	"00000001010011010110100000100000" when X"00000048",	--Add r13, r10, r13
		--	"00100001100011000000000000000001" when X"0000004c",	--Addi r12, 12, 1
		--	"00001000000000000000000000010001" when X"00000050",	--j 0x44
		--	"10101101010011010000000000000000" when X"00000054",	--sw r13,0(r10)
		--	"10001101010011110000000000000000" when X"00000058",	--lw r14,0(r10) 
		
		
			"00100000000001100000000000001001"	when X"00000000",					--ADDI R6,R0,8
			"00100000110000100000000000000000"	when X"00000004",			 		--ADDI R2,R6,0
			"00100000000010000000000000000001"	when X"00000008",					--ADDI r8, r0, 1
			"00100000110010010000000000000000"	when X"0000000c",					--ADDI R9, R6,0
			
			"00010001000000100000000000001000"	when X"00000010",					--BEQ R2,R8 Exit -- 1
			"00000000010010000001000000100010"	when X"00000014",					--Sub R2 R2 1
			"00100000000000110000000000000001"	when X"00000018",					--ADDI R3,R0,1
			"00100001001001100000000000000000"	when X"0000001c",					--ADDI R6,R9,0
			
			"00010000011000100000000000000011"	when X"00000020",					--BEQ R3, R2  --2
			"00000001001001100100100000100000"	when X"00000024",					--ADD R9,R9,R6
			"00100000011000110000000000000001"	when X"00000028",					--ADDI R3,R3,1
			"00001000000000000000000000001000"	when X"0000002c",					--J -- 2
			"00001000000000000000000000000100"	when X"00000030",					--J -- 1
			
			"10101100000010010000000000000010"	when X"00000034",					--sw r9,2(r0)
			"10001100000000010000000000000010"  when X"00000038",					--lw r1,2(r0)


	
		
		
		
         "00100000000000000000000000000000" when others; --nop (addi r0,r0,0)
                            
end behav;